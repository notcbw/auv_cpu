`ifndef _AUV_PKG_SV
`define _AUV_PKG_SV

package auv_pkg;

    typedef enum logic { OP1_RS1, OP1_PC } sel_op1_t;
    typedef enum logic { OP2_RS2, OP2_IMM } sel_op2_t;

endpackage

`endif
